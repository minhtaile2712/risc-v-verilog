module add4 (din, dout);
input [31:0] din;
output [31:0] dout;

assign dout = din + 4;
endmodule
